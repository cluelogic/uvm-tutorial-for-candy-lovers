//
// no_source_code.sv
//

module top;
   initial begin
      $display( "=====================================================" );
      $display( "No source code is available for Tutorial #", `TUTORIAL );
      $display( "Try another Tutorial Number"                           );
      $display( "=====================================================" );
   end
endmodule: top